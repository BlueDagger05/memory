package memory_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "pkt.sv"
        `include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "scoreboard.sv"
	`include "coverage.sv"
	`include "base_sequence.sv"
	`include "write_sequence.sv"
endpackage : memory_pkg
