package inclusion_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "reset_pkt_rst.sv"
	`include "sequencer_rst.sv"
	`include "driver_rst.sv"
	`include "monitor_rst.sv"
	`include "agent_rst.sv"
        `include "base_sequence_rst.sv"
endpackage : inclusion_pkg
