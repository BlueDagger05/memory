package inclusion_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "reset_pkt.sv"
	`include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
        `include "base_sequence.sv"
endpackage : inclusion_pkg
