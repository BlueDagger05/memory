interface reset_interface(input bit clk, reset_n);
endinterface: reset_interface

